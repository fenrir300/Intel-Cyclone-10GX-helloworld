module led_counter (
		input  wire        clock, //  counter_input.clock
		output wire [31:0] q      // counter_output.q
	);
endmodule

